library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity gold_rom is
port(
row_addr, col_addr : in std_logic_vector(3 downto 0);
dout : out std_logic_vector(7 downto 0));
end gold_rom;
architecture rtl of gold_rom is
type ram_type is array (0 to 15, 0 to 15) of
std_logic_vector(7 downto 0);
signal program: ram_type := (
    ("00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000010", "00000010", "00000100", "00000001","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000101", "00000000", "00000010", "00000011","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101"),
    ("00000000", "00000110", "00000001", "00000010","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101","00000001", "00000011", "00000001", "00000101")

    );
begin
dout <= program(conv_integer(unsigned(row_addr)), conv_integer(unsigned(col_addr)));
end rtl;